library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity acil_durdurma_asiri_yuk is
end acil_durdurma_asiri_yuk;

architecture Behavioral of acil_durdurma_asiri_yuk is

    -- DUT sinyalleri
    signal clk           : std_logic := '0';
    signal reset_n       : std_logic := '0';
    signal call_btn      : std_logic_vector(3 downto 0) := (others => '0');
    signal cab_btn       : std_logic_vector(3 downto 0) := (others => '0');
    signal overload      : std_logic := '0';
    signal emergency     : std_logic := '0';

    signal current_floor : std_logic_vector(1 downto 0);
    signal motor_up      : std_logic;
    signal motor_down    : std_logic;
    signal door_open     : std_logic;
    signal door_close    : std_logic;

    constant CLK_PERIOD : time := 10 ns;

begin

    ----------------------------------------------------------------
    -- DUT bağlama
    ----------------------------------------------------------------
    DUT: entity work.main
        port map (
            clk           => clk,
            reset_n       => reset_n,
            call_btn      => call_btn,
            cab_btn       => cab_btn,
            overload      => overload,
            emergency     => emergency,
            current_floor => current_floor,
            motor_up      => motor_up,
            motor_down    => motor_down,
            door_open     => door_open,
            door_close    => door_close
        );

    ----------------------------------------------------------------
    -- Clock üretimi
    ----------------------------------------------------------------
    clk_process : process
    begin
        while true loop
            clk <= '0';
            wait for CLK_PERIOD/2;
            clk <= '1';
            wait for CLK_PERIOD/2;
        end loop;
    end process;

    ----------------------------------------------------------------
    -- Test senaryosu
    ----------------------------------------------------------------
    stim_proc: process
    begin
        -- Reset
        reset_n <= '0';
        wait for 50 ns;
        reset_n <= '1';

        -- Kat 2 çağrısı (kapı açma ve motor hareket test)
        call_btn(2) <= '1';
        wait for 20 ns;
        call_btn(2) <= '0';

        -- Asansör kat 2'ye doğru hareket ederken overload testi
        wait for 100 ns;
        overload <= '1'; -- overload geldi, kapı açık kalmalı
        wait for 50 ns;
        overload <= '0'; -- overload kalktı, kapı kapanabilir

        -- Kabin içi çağrı testi
        cab_btn(0) <= '1';
        wait for 20 ns;
        cab_btn(0) <= '0';

        -- Acil durum testi
        wait for 100 ns;
        emergency <= '1'; -- acil durum, kapı açık kalmalı
        wait for 50 ns;
        emergency <= '0';

        -- Simülasyon bitiş
        wait for 200 ns;
        assert false report "Simulation ended" severity note;
        wait;
    end process;

end Behavioral;
